/****************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            ARPS_IP_master_seq_lib.sv

    DESCRIPTION     sequence includes

 ****************************************************************************/

`ifndef ARPS_IP_AXIL_SEQ_LIB_SV
`define ARPS_IP_AXIL_SEQ_LIB_SV

`include "sequences/ARPS_IP_axil_base_seq.sv"
`include "sequences/ARPS_IP_axil_simple_seq.sv"

`endif
