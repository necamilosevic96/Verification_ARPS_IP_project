library verilog;
use verilog.vl_types.all;
entity ARPS_IP_pkg_sv_unit is
end ARPS_IP_pkg_sv_unit;
