/****************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            ARPS_IP_test_lib.sv

    DESCRIPTION     test includes

 ****************************************************************************/

`ifndef ARPS_IP_TEST_LIB_SV
`define ARPS_IP_TEST_LIB_SV

`include "ARPS_IP_test_base.sv"
`include "ARPS_IP_test_simple.sv"
    
`endif
