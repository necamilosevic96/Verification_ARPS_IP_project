library verilog;
use verilog.vl_types.all;
entity axil_if is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end axil_if;
