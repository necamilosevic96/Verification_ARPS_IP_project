library verilog;
use verilog.vl_types.all;
entity ARPS_IP_test_top is
end ARPS_IP_test_top;
