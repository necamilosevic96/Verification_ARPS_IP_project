/****************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            ARPS_IP_master_seq_lib.sv

    DESCRIPTION     sequence includes

 ****************************************************************************/

`ifndef ARPS_IP_BRAM_CURR_SEQ_LIB_SV
`define ARPS_IP_BRAM_CURR_SEQ_LIB_SV

`include "sequences/ARPS_IP_bram_curr_base_seq.sv"
`include "sequences/ARPS_IP_bram_curr_simple_seq.sv"
`include "sequences/ARPS_IP_bram_curr_base_seq_2.sv"
`include "sequences/ARPS_IP_bram_curr_simple_seq_2.sv"

`endif
