library verilog;
use verilog.vl_types.all;
entity ARPS_IP_pkg is
end ARPS_IP_pkg;
